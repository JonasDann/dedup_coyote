    // ----------------------------------------------------------------------
    // USER 
    // ----------------------------------------------------------------------
    dedup_4k inst_dedup ( 
        .axi_ctrl_araddr        (axi_ctrl.araddr[16-1:0]), // use LSBs (high-bits start with 0x8xxx)
        .axi_ctrl_arprot        (axi_ctrl.arprot),
        .axi_ctrl_arready       (axi_ctrl.arready),
        .axi_ctrl_arvalid       (axi_ctrl.arvalid),
        .axi_ctrl_awaddr        (axi_ctrl.awaddr[16-1:0]),
        .axi_ctrl_awprot        (axi_ctrl.awprot),
        .axi_ctrl_awready       (axi_ctrl.awready),
        .axi_ctrl_awvalid       (axi_ctrl.awvalid),
        .axi_ctrl_bready        (axi_ctrl.bready),
        .axi_ctrl_bresp         (axi_ctrl.bresp),
        .axi_ctrl_bvalid        (axi_ctrl.bvalid),
        .axi_ctrl_rdata         (axi_ctrl.rdata),
        .axi_ctrl_rready        (axi_ctrl.rready),
        .axi_ctrl_rresp         (axi_ctrl.rresp),
        .axi_ctrl_rvalid        (axi_ctrl.rvalid),
        .axi_ctrl_wdata         (axi_ctrl.wdata),
        .axi_ctrl_wready        (axi_ctrl.wready),
        .axi_ctrl_wstrb         (axi_ctrl.wstrb),
        .axi_ctrl_wvalid        (axi_ctrl.wvalid),

        .hostd_bpss_rd_req_valid      (bpss_rd_req.valid),
        .hostd_bpss_rd_req_ready      (bpss_rd_req.ready),
        .hostd_bpss_rd_req_data       (bpss_rd_req.data),
        .hostd_bpss_wr_req_valid      (bpss_wr_req.valid),
        .hostd_bpss_wr_req_ready      (bpss_wr_req.ready),
        .hostd_bpss_wr_req_data       (bpss_wr_req.data),
        .hostd_bpss_rd_done_valid     (bpss_rd_done.valid),
        .hostd_bpss_rd_done_ready     (bpss_rd_done.ready),
        .hostd_bpss_rd_done_data      (bpss_rd_done.data),
        .hostd_bpss_wr_done_valid     (bpss_wr_done.valid),
        .hostd_bpss_wr_done_ready     (bpss_wr_done.ready),
        .hostd_bpss_wr_done_data      (bpss_wr_done.data),
        .hostd_axis_host_sink_tdata   (axis_host_0_sink.tdata),
        .hostd_axis_host_sink_tkeep   (axis_host_0_sink.tkeep),
        .hostd_axis_host_sink_tlast   (axis_host_0_sink.tlast),
        .hostd_axis_host_sink_tready  (axis_host_0_sink.tready),
        .hostd_axis_host_sink_tvalid  (axis_host_0_sink.tvalid),
        .hostd_axis_host_src_tdata    (axis_host_0_src.tdata),
        .hostd_axis_host_src_tkeep    (axis_host_0_src.tkeep),
        .hostd_axis_host_src_tlast    (axis_host_0_src.tlast),
        .hostd_axis_host_src_tready   (axis_host_0_src.tready),
        .hostd_axis_host_src_tvalid   (axis_host_0_src.tvalid),

        .networkIo_rdma_0_sq_valid           (rdma_0_sq.valid         ),
        .networkIo_rdma_0_sq_ready           (rdma_0_sq.ready         ),
        .networkIo_rdma_0_sq_data            (rdma_0_sq.data          ),
        .networkIo_rdma_0_ack_valid          (rdma_0_ack.valid        ),
        .networkIo_rdma_0_ack_ready          (rdma_0_ack.ready        ),
        .networkIo_rdma_0_ack_data           (rdma_0_ack.data         ),
        .networkIo_rdma_0_rd_req_valid       (rdma_0_rd_req.valid     ),
        .networkIo_rdma_0_rd_req_ready       (rdma_0_rd_req.ready     ),
        .networkIo_rdma_0_rd_req_data        (rdma_0_rd_req.data      ),
        .networkIo_rdma_0_wr_req_valid       (rdma_0_wr_req.valid     ),
        .networkIo_rdma_0_wr_req_ready       (rdma_0_wr_req.ready     ),
        .networkIo_rdma_0_wr_req_data        (rdma_0_wr_req.data      ),
        .networkIo_axis_rdma_0_sink_tvalid   (axis_rdma_0_sink.tvalid ),
        .networkIo_axis_rdma_0_sink_tready   (axis_rdma_0_sink.tready ),
        .networkIo_axis_rdma_0_sink_tdata    (axis_rdma_0_sink.tdata  ),
        .networkIo_axis_rdma_0_sink_tkeep    (axis_rdma_0_sink.tkeep  ),
        .networkIo_axis_rdma_0_sink_tid      (axis_rdma_0_sink.tid    ),
        .networkIo_axis_rdma_0_sink_tlast    (axis_rdma_0_sink.tlast  ),
        .networkIo_axis_rdma_0_src_tvalid    (axis_rdma_0_src.tvalid  ),
        .networkIo_axis_rdma_0_src_tready    (axis_rdma_0_src.tready  ),
        .networkIo_axis_rdma_0_src_tdata     (axis_rdma_0_src.tdata   ),
        .networkIo_axis_rdma_0_src_tkeep     (axis_rdma_0_src.tkeep   ),
        .networkIo_axis_rdma_0_src_tid       (axis_rdma_0_src.tid     ),
        .networkIo_axis_rdma_0_src_tlast     (axis_rdma_0_src.tlast   ),
        .axi_mem_0_araddr(axi_mem_0_araddr),
        .axi_mem_0_arburst(axi_mem_0_arburst),
        //.axi_mem_0_arcache(axi_mem_0_arcache),
        .axi_mem_0_arid(axi_mem_0_arid),
        .axi_mem_0_arlen(axi_mem_0_arlen),
        //.axi_mem_0_arlock(axi_mem_0_arlock),
        //.axi_mem_0_arprot(axi_mem_0_arprot),
        //.axi_mem_0_arqos(axi_mem_0_arqos),
        .axi_mem_0_arready(axi_mem_0_arready),
        //.axi_mem_0_arregion(axi_mem_0_arregion),
        .axi_mem_0_arsize(axi_mem_0_arsize),
        .axi_mem_0_arvalid(axi_mem_0_arvalid),
        .axi_mem_0_awaddr(axi_mem_0_awaddr),
        .axi_mem_0_awburst(axi_mem_0_awburst),
        //.axi_mem_0_awcache(axi_mem_0_awcache),
        .axi_mem_0_awid(axi_mem_0_awid),
        .axi_mem_0_awlen(axi_mem_0_awlen),
        //.axi_mem_0_awlock(axi_mem_0_awlock),
        //.axi_mem_0_awprot(axi_mem_0_awprot),
        //.axi_mem_0_awqos(axi_mem_0_awqos),
        .axi_mem_0_awready(axi_mem_0_awready),
        //.axi_mem_0_awregion(axi_mem_0_awregion),
        .axi_mem_0_awsize(axi_mem_0_awsize),
        .axi_mem_0_awvalid(axi_mem_0_awvalid),
        .axi_mem_0_bid(axi_mem_0_bid),
        .axi_mem_0_bready(axi_mem_0_bready),
        .axi_mem_0_bresp(axi_mem_0_bresp),
        .axi_mem_0_bvalid(axi_mem_0_bvalid),
        .axi_mem_0_rdata(axi_mem_0_rdata),
        .axi_mem_0_rid(axi_mem_0_rid),
        .axi_mem_0_rlast(axi_mem_0_rlast),
        .axi_mem_0_rready(axi_mem_0_rready),
        .axi_mem_0_rresp(axi_mem_0_rresp),
        .axi_mem_0_rvalid(axi_mem_0_rvalid),
        .axi_mem_0_wdata(axi_mem_0_wdata),
        .axi_mem_0_wlast(axi_mem_0_wlast),
        .axi_mem_0_wready(axi_mem_0_wready),
        .axi_mem_0_wstrb(axi_mem_0_wstrb),
        .axi_mem_0_wvalid(axi_mem_0_wvalid),
        .axi_mem_1_araddr(axi_mem_1_araddr),
        .axi_mem_1_arburst(axi_mem_1_arburst),
        //.axi_mem_1_arcache(axi_mem_1_arcache),
        .axi_mem_1_arid(axi_mem_1_arid),
        .axi_mem_1_arlen(axi_mem_1_arlen),
        //.axi_mem_1_arlock(axi_mem_1_arlock),
        //.axi_mem_1_arprot(axi_mem_1_arprot),
        //.axi_mem_1_arqos(axi_mem_1_arqos),
        .axi_mem_1_arready(axi_mem_1_arready),
        //.axi_mem_1_arregion(axi_mem_1_arregion),
        .axi_mem_1_arsize(axi_mem_1_arsize),
        .axi_mem_1_arvalid(axi_mem_1_arvalid),
        .axi_mem_1_awaddr(axi_mem_1_awaddr),
        .axi_mem_1_awburst(axi_mem_1_awburst),
        //.axi_mem_1_awcache(axi_mem_1_awcache),
        .axi_mem_1_awid(axi_mem_1_awid),
        .axi_mem_1_awlen(axi_mem_1_awlen),
        //.axi_mem_1_awlock(axi_mem_1_awlock),
        //.axi_mem_1_awprot(axi_mem_1_awprot),
        //.axi_mem_1_awqos(axi_mem_1_awqos),
        .axi_mem_1_awready(axi_mem_1_awready),
        //.axi_mem_1_awregion(axi_mem_1_awregion),
        .axi_mem_1_awsize(axi_mem_1_awsize),
        .axi_mem_1_awvalid(axi_mem_1_awvalid),
        .axi_mem_1_bid(axi_mem_1_bid),
        .axi_mem_1_bready(axi_mem_1_bready),
        .axi_mem_1_bresp(axi_mem_1_bresp),
        .axi_mem_1_bvalid(axi_mem_1_bvalid),
        .axi_mem_1_rdata(axi_mem_1_rdata),
        .axi_mem_1_rid(axi_mem_1_rid),
        .axi_mem_1_rlast(axi_mem_1_rlast),
        .axi_mem_1_rready(axi_mem_1_rready),
        .axi_mem_1_rresp(axi_mem_1_rresp),
        .axi_mem_1_rvalid(axi_mem_1_rvalid),
        .axi_mem_1_wdata(axi_mem_1_wdata),
        .axi_mem_1_wlast(axi_mem_1_wlast),
        .axi_mem_1_wready(axi_mem_1_wready),
        .axi_mem_1_wstrb(axi_mem_1_wstrb),
        .axi_mem_1_wvalid(axi_mem_1_wvalid),
        .axi_mem_2_araddr(axi_mem_2_araddr),
        .axi_mem_2_arburst(axi_mem_2_arburst),
        //.axi_mem_2_arcache(axi_mem_2_arcache),
        .axi_mem_2_arid(axi_mem_2_arid),
        .axi_mem_2_arlen(axi_mem_2_arlen),
        //.axi_mem_2_arlock(axi_mem_2_arlock),
        //.axi_mem_2_arprot(axi_mem_2_arprot),
        //.axi_mem_2_arqos(axi_mem_2_arqos),
        .axi_mem_2_arready(axi_mem_2_arready),
        //.axi_mem_2_arregion(axi_mem_2_arregion),
        .axi_mem_2_arsize(axi_mem_2_arsize),
        .axi_mem_2_arvalid(axi_mem_2_arvalid),
        .axi_mem_2_awaddr(axi_mem_2_awaddr),
        .axi_mem_2_awburst(axi_mem_2_awburst),
        //.axi_mem_2_awcache(axi_mem_2_awcache),
        .axi_mem_2_awid(axi_mem_2_awid),
        .axi_mem_2_awlen(axi_mem_2_awlen),
        //.axi_mem_2_awlock(axi_mem_2_awlock),
        //.axi_mem_2_awprot(axi_mem_2_awprot),
        //.axi_mem_2_awqos(axi_mem_2_awqos),
        .axi_mem_2_awready(axi_mem_2_awready),
        //.axi_mem_2_awregion(axi_mem_2_awregion),
        .axi_mem_2_awsize(axi_mem_2_awsize),
        .axi_mem_2_awvalid(axi_mem_2_awvalid),
        .axi_mem_2_bid(axi_mem_2_bid),
        .axi_mem_2_bready(axi_mem_2_bready),
        .axi_mem_2_bresp(axi_mem_2_bresp),
        .axi_mem_2_bvalid(axi_mem_2_bvalid),
        .axi_mem_2_rdata(axi_mem_2_rdata),
        .axi_mem_2_rid(axi_mem_2_rid),
        .axi_mem_2_rlast(axi_mem_2_rlast),
        .axi_mem_2_rready(axi_mem_2_rready),
        .axi_mem_2_rresp(axi_mem_2_rresp),
        .axi_mem_2_rvalid(axi_mem_2_rvalid),
        .axi_mem_2_wdata(axi_mem_2_wdata),
        .axi_mem_2_wlast(axi_mem_2_wlast),
        .axi_mem_2_wready(axi_mem_2_wready),
        .axi_mem_2_wstrb(axi_mem_2_wstrb),
        .axi_mem_2_wvalid(axi_mem_2_wvalid),
        .axi_mem_3_araddr(axi_mem_3_araddr),
        .axi_mem_3_arburst(axi_mem_3_arburst),
        //.axi_mem_3_arcache(axi_mem_3_arcache),
        .axi_mem_3_arid(axi_mem_3_arid),
        .axi_mem_3_arlen(axi_mem_3_arlen),
        //.axi_mem_3_arlock(axi_mem_3_arlock),
        //.axi_mem_3_arprot(axi_mem_3_arprot),
        //.axi_mem_3_arqos(axi_mem_3_arqos),
        .axi_mem_3_arready(axi_mem_3_arready),
        //.axi_mem_3_arregion(axi_mem_3_arregion),
        .axi_mem_3_arsize(axi_mem_3_arsize),
        .axi_mem_3_arvalid(axi_mem_3_arvalid),
        .axi_mem_3_awaddr(axi_mem_3_awaddr),
        .axi_mem_3_awburst(axi_mem_3_awburst),
        //.axi_mem_3_awcache(axi_mem_3_awcache),
        .axi_mem_3_awid(axi_mem_3_awid),
        .axi_mem_3_awlen(axi_mem_3_awlen),
        //.axi_mem_3_awlock(axi_mem_3_awlock),
        //.axi_mem_3_awprot(axi_mem_3_awprot),
        //.axi_mem_3_awqos(axi_mem_3_awqos),
        .axi_mem_3_awready(axi_mem_3_awready),
        //.axi_mem_3_awregion(axi_mem_3_awregion),
        .axi_mem_3_awsize(axi_mem_3_awsize),
        .axi_mem_3_awvalid(axi_mem_3_awvalid),
        .axi_mem_3_bid(axi_mem_3_bid),
        .axi_mem_3_bready(axi_mem_3_bready),
        .axi_mem_3_bresp(axi_mem_3_bresp),
        .axi_mem_3_bvalid(axi_mem_3_bvalid),
        .axi_mem_3_rdata(axi_mem_3_rdata),
        .axi_mem_3_rid(axi_mem_3_rid),
        .axi_mem_3_rlast(axi_mem_3_rlast),
        .axi_mem_3_rready(axi_mem_3_rready),
        .axi_mem_3_rresp(axi_mem_3_rresp),
        .axi_mem_3_rvalid(axi_mem_3_rvalid),
        .axi_mem_3_wdata(axi_mem_3_wdata),
        .axi_mem_3_wlast(axi_mem_3_wlast),
        .axi_mem_3_wready(axi_mem_3_wready),
        .axi_mem_3_wstrb(axi_mem_3_wstrb),
        .axi_mem_3_wvalid(axi_mem_3_wvalid),
        .axi_mem_4_araddr(axi_mem_4_araddr),
        .axi_mem_4_arburst(axi_mem_4_arburst),
        //.axi_mem_4_arcache(axi_mem_4_arcache),
        .axi_mem_4_arid(axi_mem_4_arid),
        .axi_mem_4_arlen(axi_mem_4_arlen),
        //.axi_mem_4_arlock(axi_mem_4_arlock),
        //.axi_mem_4_arprot(axi_mem_4_arprot),
        //.axi_mem_4_arqos(axi_mem_4_arqos),
        .axi_mem_4_arready(axi_mem_4_arready),
        //.axi_mem_4_arregion(axi_mem_4_arregion),
        .axi_mem_4_arsize(axi_mem_4_arsize),
        .axi_mem_4_arvalid(axi_mem_4_arvalid),
        .axi_mem_4_awaddr(axi_mem_4_awaddr),
        .axi_mem_4_awburst(axi_mem_4_awburst),
        //.axi_mem_4_awcache(axi_mem_4_awcache),
        .axi_mem_4_awid(axi_mem_4_awid),
        .axi_mem_4_awlen(axi_mem_4_awlen),
        //.axi_mem_4_awlock(axi_mem_4_awlock),
        //.axi_mem_4_awprot(axi_mem_4_awprot),
        //.axi_mem_4_awqos(axi_mem_4_awqos),
        .axi_mem_4_awready(axi_mem_4_awready),
        //.axi_mem_4_awregion(axi_mem_4_awregion),
        .axi_mem_4_awsize(axi_mem_4_awsize),
        .axi_mem_4_awvalid(axi_mem_4_awvalid),
        .axi_mem_4_bid(axi_mem_4_bid),
        .axi_mem_4_bready(axi_mem_4_bready),
        .axi_mem_4_bresp(axi_mem_4_bresp),
        .axi_mem_4_bvalid(axi_mem_4_bvalid),
        .axi_mem_4_rdata(axi_mem_4_rdata),
        .axi_mem_4_rid(axi_mem_4_rid),
        .axi_mem_4_rlast(axi_mem_4_rlast),
        .axi_mem_4_rready(axi_mem_4_rready),
        .axi_mem_4_rresp(axi_mem_4_rresp),
        .axi_mem_4_rvalid(axi_mem_4_rvalid),
        .axi_mem_4_wdata(axi_mem_4_wdata),
        .axi_mem_4_wlast(axi_mem_4_wlast),
        .axi_mem_4_wready(axi_mem_4_wready),
        .axi_mem_4_wstrb(axi_mem_4_wstrb),
        .axi_mem_4_wvalid(axi_mem_4_wvalid),

        .axi_mem_5_araddr(axi_mem_5_araddr),
        .axi_mem_5_arburst(axi_mem_5_arburst),
        //.axi_mem_5_arcache(axi_mem_5_arcache),
        .axi_mem_5_arid(axi_mem_5_arid),
        .axi_mem_5_arlen(axi_mem_5_arlen),
        //.axi_mem_5_arlock(axi_mem_5_arlock),
        //.axi_mem_5_arprot(axi_mem_5_arprot),
        //.axi_mem_5_arqos(axi_mem_5_arqos),
        .axi_mem_5_arready(axi_mem_5_arready),
        //.axi_mem_5_arregion(axi_mem_5_arregion),
        .axi_mem_5_arsize(axi_mem_5_arsize),
        .axi_mem_5_arvalid(axi_mem_5_arvalid),
        .axi_mem_5_awaddr(axi_mem_5_awaddr),
        .axi_mem_5_awburst(axi_mem_5_awburst),
        //.axi_mem_5_awcache(axi_mem_5_awcache),
        .axi_mem_5_awid(axi_mem_5_awid),
        .axi_mem_5_awlen(axi_mem_5_awlen),
        //.axi_mem_5_awlock(axi_mem_5_awlock),
        //.axi_mem_5_awprot(axi_mem_5_awprot),
        //.axi_mem_5_awqos(axi_mem_5_awqos),
        .axi_mem_5_awready(axi_mem_5_awready),
        //.axi_mem_5_awregion(axi_mem_5_awregion),
        .axi_mem_5_awsize(axi_mem_5_awsize),
        .axi_mem_5_awvalid(axi_mem_5_awvalid),
        .axi_mem_5_bid(axi_mem_5_bid),
        .axi_mem_5_bready(axi_mem_5_bready),
        .axi_mem_5_bresp(axi_mem_5_bresp),
        .axi_mem_5_bvalid(axi_mem_5_bvalid),
        .axi_mem_5_rdata(axi_mem_5_rdata),
        .axi_mem_5_rid(axi_mem_5_rid),
        .axi_mem_5_rlast(axi_mem_5_rlast),
        .axi_mem_5_rready(axi_mem_5_rready),
        .axi_mem_5_rresp(axi_mem_5_rresp),
        .axi_mem_5_rvalid(axi_mem_5_rvalid),
        .axi_mem_5_wdata(axi_mem_5_wdata),
        .axi_mem_5_wlast(axi_mem_5_wlast),
        .axi_mem_5_wready(axi_mem_5_wready),
        .axi_mem_5_wstrb(axi_mem_5_wstrb),
        .axi_mem_5_wvalid(axi_mem_5_wvalid),

        .axi_mem_6_araddr(axi_mem_6_araddr),
        .axi_mem_6_arburst(axi_mem_6_arburst),
        //.axi_mem_6_arcache(axi_mem_6_arcache),
        .axi_mem_6_arid(axi_mem_6_arid),
        .axi_mem_6_arlen(axi_mem_6_arlen),
        //.axi_mem_6_arlock(axi_mem_6_arlock),
        //.axi_mem_6_arprot(axi_mem_6_arprot),
        //.axi_mem_6_arqos(axi_mem_6_arqos),
        .axi_mem_6_arready(axi_mem_6_arready),
        //.axi_mem_6_arregion(axi_mem_6_arregion),
        .axi_mem_6_arsize(axi_mem_6_arsize),
        .axi_mem_6_arvalid(axi_mem_6_arvalid),
        .axi_mem_6_awaddr(axi_mem_6_awaddr),
        .axi_mem_6_awburst(axi_mem_6_awburst),
        //.axi_mem_6_awcache(axi_mem_6_awcache),
        .axi_mem_6_awid(axi_mem_6_awid),
        .axi_mem_6_awlen(axi_mem_6_awlen),
        //.axi_mem_6_awlock(axi_mem_6_awlock),
        //.axi_mem_6_awprot(axi_mem_6_awprot),
        //.axi_mem_6_awqos(axi_mem_6_awqos),
        .axi_mem_6_awready(axi_mem_6_awready),
        //.axi_mem_6_awregion(axi_mem_6_awregion),
        .axi_mem_6_awsize(axi_mem_6_awsize),
        .axi_mem_6_awvalid(axi_mem_6_awvalid),
        .axi_mem_6_bid(axi_mem_6_bid),
        .axi_mem_6_bready(axi_mem_6_bready),
        .axi_mem_6_bresp(axi_mem_6_bresp),
        .axi_mem_6_bvalid(axi_mem_6_bvalid),
        .axi_mem_6_rdata(axi_mem_6_rdata),
        .axi_mem_6_rid(axi_mem_6_rid),
        .axi_mem_6_rlast(axi_mem_6_rlast),
        .axi_mem_6_rready(axi_mem_6_rready),
        .axi_mem_6_rresp(axi_mem_6_rresp),
        .axi_mem_6_rvalid(axi_mem_6_rvalid),
        .axi_mem_6_wdata(axi_mem_6_wdata),
        .axi_mem_6_wlast(axi_mem_6_wlast),
        .axi_mem_6_wready(axi_mem_6_wready),
        .axi_mem_6_wstrb(axi_mem_6_wstrb),
        .axi_mem_6_wvalid(axi_mem_6_wvalid),

        // .axi_mem_7_araddr(axi_mem_7_araddr),
        // .axi_mem_7_arburst(axi_mem_7_arburst),
        // //.axi_mem_7_arcache(axi_mem_7_arcache),
        // .axi_mem_7_arid(axi_mem_7_arid),
        // .axi_mem_7_arlen(axi_mem_7_arlen),
        // //.axi_mem_7_arlock(axi_mem_7_arlock),
        // //.axi_mem_7_arprot(axi_mem_7_arprot),
        // //.axi_mem_7_arqos(axi_mem_7_arqos),
        // .axi_mem_7_arready(axi_mem_7_arready),
        // //.axi_mem_7_arregion(axi_mem_7_arregion),
        // .axi_mem_7_arsize(axi_mem_7_arsize),
        // .axi_mem_7_arvalid(axi_mem_7_arvalid),
        // .axi_mem_7_awaddr(axi_mem_7_awaddr),
        // .axi_mem_7_awburst(axi_mem_7_awburst),
        // //.axi_mem_7_awcache(axi_mem_7_awcache),
        // .axi_mem_7_awid(axi_mem_7_awid),
        // .axi_mem_7_awlen(axi_mem_7_awlen),
        // //.axi_mem_7_awlock(axi_mem_7_awlock),
        // //.axi_mem_7_awprot(axi_mem_7_awprot),
        // //.axi_mem_7_awqos(axi_mem_7_awqos),
        // .axi_mem_7_awready(axi_mem_7_awready),
        // //.axi_mem_7_awregion(axi_mem_7_awregion),
        // .axi_mem_7_awsize(axi_mem_7_awsize),
        // .axi_mem_7_awvalid(axi_mem_7_awvalid),
        // .axi_mem_7_bid(axi_mem_7_bid),
        // .axi_mem_7_bready(axi_mem_7_bready),
        // .axi_mem_7_bresp(axi_mem_7_bresp),
        // .axi_mem_7_bvalid(axi_mem_7_bvalid),
        // .axi_mem_7_rdata(axi_mem_7_rdata),
        // .axi_mem_7_rid(axi_mem_7_rid),
        // .axi_mem_7_rlast(axi_mem_7_rlast),
        // .axi_mem_7_rready(axi_mem_7_rready),
        // .axi_mem_7_rresp(axi_mem_7_rresp),
        // .axi_mem_7_rvalid(axi_mem_7_rvalid),
        // .axi_mem_7_wdata(axi_mem_7_wdata),
        // .axi_mem_7_wlast(axi_mem_7_wlast),
        // .axi_mem_7_wready(axi_mem_7_wready),
        // .axi_mem_7_wstrb(axi_mem_7_wstrb),
        // .axi_mem_7_wvalid(axi_mem_7_wvalid),

        // .axi_mem_8_araddr(axi_mem_8_araddr),
        // .axi_mem_8_arburst(axi_mem_8_arburst),
        // //.axi_mem_8_arcache(axi_mem_8_arcache),
        // .axi_mem_8_arid(axi_mem_8_arid),
        // .axi_mem_8_arlen(axi_mem_8_arlen),
        // //.axi_mem_8_arlock(axi_mem_8_arlock),
        // //.axi_mem_8_arprot(axi_mem_8_arprot),
        // //.axi_mem_8_arqos(axi_mem_8_arqos),
        // .axi_mem_8_arready(axi_mem_8_arready),
        // //.axi_mem_8_arregion(axi_mem_8_arregion),
        // .axi_mem_8_arsize(axi_mem_8_arsize),
        // .axi_mem_8_arvalid(axi_mem_8_arvalid),
        // .axi_mem_8_awaddr(axi_mem_8_awaddr),
        // .axi_mem_8_awburst(axi_mem_8_awburst),
        // //.axi_mem_8_awcache(axi_mem_8_awcache),
        // .axi_mem_8_awid(axi_mem_8_awid),
        // .axi_mem_8_awlen(axi_mem_8_awlen),
        // //.axi_mem_8_awlock(axi_mem_8_awlock),
        // //.axi_mem_8_awprot(axi_mem_8_awprot),
        // //.axi_mem_8_awqos(axi_mem_8_awqos),
        // .axi_mem_8_awready(axi_mem_8_awready),
        // //.axi_mem_8_awregion(axi_mem_8_awregion),
        // .axi_mem_8_awsize(axi_mem_8_awsize),
        // .axi_mem_8_awvalid(axi_mem_8_awvalid),
        // .axi_mem_8_bid(axi_mem_8_bid),
        // .axi_mem_8_bready(axi_mem_8_bready),
        // .axi_mem_8_bresp(axi_mem_8_bresp),
        // .axi_mem_8_bvalid(axi_mem_8_bvalid),
        // .axi_mem_8_rdata(axi_mem_8_rdata),
        // .axi_mem_8_rid(axi_mem_8_rid),
        // .axi_mem_8_rlast(axi_mem_8_rlast),
        // .axi_mem_8_rready(axi_mem_8_rready),
        // .axi_mem_8_rresp(axi_mem_8_rresp),
        // .axi_mem_8_rvalid(axi_mem_8_rvalid),
        // .axi_mem_8_wdata(axi_mem_8_wdata),
        // .axi_mem_8_wlast(axi_mem_8_wlast),
        // .axi_mem_8_wready(axi_mem_8_wready),
        // .axi_mem_8_wstrb(axi_mem_8_wstrb),
        // .axi_mem_8_wvalid(axi_mem_8_wvalid),

        .clk                   (aclk),
        .resetn                (aresetn)
    );